library verilog;
use verilog.vl_types.all;
entity Morse_vlg_vec_tst is
end Morse_vlg_vec_tst;
