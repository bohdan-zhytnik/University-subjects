library verilog;
use verilog.vl_types.all;
entity MorseZHYT_vlg_vec_tst is
end MorseZHYT_vlg_vec_tst;
