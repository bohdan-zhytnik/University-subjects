-- Character ROM font Consolas 24 pts from 32 to 127 ASCII character
-- Charter size width = 24, height 32;
-- The file has the structure that compiles exactly to 9 memory M9K blocks. 
library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all;

entity Consolas24pt_Font is
	port(clk: in std_logic;
		addr: in std_logic_vector(11 downto 0);
		fontRow: out std_logic_vector(0 to 23)
	);
end entity;

architecture Behavioral of Consolas24pt_Font is
 
	type rom_type is array (0 to 3071) of std_logic_vector(0 to 23);
	-- ROM definition
	signal ROM : rom_type := (   
-- char code 32 0x20 Space
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  --  
 X"000000",   --  
-- char code 33 0x21 Exclamation mark
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"000000", -- 
 X"000000", -- 
 X"00c000", --          ##
 X"01e000", --         ####
 X"01e000", --         ####
 X"00c000", --          ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 34 0x22 Quotation mark
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"0f1e00", --      ####   ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 35 0x23 Number sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"031c00", --        ##   ###
 X"031c00", --        ##   ###
 X"031c00", --        ##   ###
 X"031c00", --        ##   ###
 X"031c00", --        ##   ###
 X"3fff80", --    ###############
 X"3fff80", --    ###############
 X"073800", --       ###  ###
 X"073800", --       ###  ###
 X"073800", --       ###  ###
 X"063800", --       ##   ###
 X"063800", --       ##   ###
 X"7fff00", --   ###############
 X"7fff00", --   ###############
 X"063800", --       ##   ###
 X"0e7000", --      ###  ###
 X"0e7000", --      ###  ###
 X"0e7000", --      ###  ###
 X"0e7000", --      ###  ###
 X"0e7000", --      ###  ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 36 0x24 Dollar sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"003000", --            ##
 X"003000", --            ##
 X"007000", --           ###
 X"03fc00", --        ########
 X"0ffe00", --      ###########
 X"1e6200", --     ####  ##   #
 X"386000", --    ###    ##
 X"386000", --    ###    ##
 X"386000", --    ###    ##
 X"3ce000", --    ####  ###
 X"1ee000", --     #### ###
 X"1fc000", --     #######
 X"07f000", --       #######
 X"01fc00", --         #######
 X"00fe00", --          #######
 X"00cf00", --          ##  ####
 X"01c700", --         ###   ###
 X"01c700", --         ###   ###
 X"018700", --         ##    ###
 X"018f00", --         ##   ####
 X"319e00", --    ##   ##  ####
 X"3ffc00", --    ############
 X"0ff000", --      ########
 X"018000", --         ##
 X"038000", --        ###
 X"038000", --        ###
 X"030000", --        ##
 X"000000", -- 
 X"000000", -- 
-- char code 37 0x25 Percent sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1f0180", --     #####       ##
 X"3f8380", --    #######     ###
 X"79c700", --   ####  ###   ###
 X"71c600", --   ###   ###   ##
 X"71ce00", --   ###   ###  ###
 X"71dc00", --   ###   ### ###
 X"73d800", --   ###  #### ##
 X"3fb000", --    ####### ##
 X"1f7000", --     ##### ###
 X"006000", --           ##
 X"00c000", --          ##
 X"01c000", --         ###
 X"038000", --        ###
 X"031f00", --        ##   #####
 X"073f80", --       ###  #######
 X"0e79c0", --      ###  ####  ###
 X"0c71c0", --      ##   ###   ###
 X"1c71c0", --     ###   ###   ###
 X"3871c0", --    ###    ###   ###
 X"3073c0", --    ##     ###  ####
 X"703f80", --   ###      #######
 X"e01f00", --  ###        #####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 38 0x26 Ampersand
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03e000", --        #####
 X"0ff000", --      ########
 X"0e7800", --      ###  ####
 X"1c3800", --     ###    ###
 X"1c3800", --     ###    ###
 X"1c3800", --     ###    ###
 X"1c3800", --     ###    ###
 X"1e7000", --     ####  ###
 X"0fe000", --      #######
 X"0fc000", --      ######
 X"0f8000", --      #####
 X"1f8700", --     ######    ###
 X"3dc700", --    #### ###   ###
 X"38e700", --    ###   ###  ###
 X"70f700", --   ###    #### ###
 X"707e00", --   ###     ######
 X"703e00", --   ###      #####
 X"701e00", --   ###       ####
 X"781e00", --   ####      ####
 X"3c3f00", --    ####    ######
 X"1ff780", --     ######### ####
 X"0fc3c0", --      ######    ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 39 0x27 Apostrophe
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 40 0x28 Left parenthesis
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"001000", --             #
 X"003800", --            ###
 X"007000", --           ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"038000", --        ###
 X"038000", --        ###
 X"070000", --       ###
 X"070000", --       ###
 X"060000", --       ##
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0f0000", --      ####
 X"070000", --       ###
 X"070000", --       ###
 X"038000", --        ###
 X"038000", --        ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"00e000", --          ###
 X"007000", --           ###
 X"003800", --            ###
 X"001000", --             #
-- char code 41 0x29 Right parenthesis
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"040000", --       #
 X"0e0000", --      ###
 X"070000", --       ###
 X"038000", --        ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"007000", --           ###
 X"007000", --           ###
 X"007800", --           ####
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"007000", --           ###
 X"007000", --           ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"038000", --        ###
 X"070000", --       ###
 X"0e0000", --      ###
 X"040000", --       #
-- char code 42 0x2A Asterisk
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00c000", --          ##
 X"00c000", --          ##
 X"08c400", --      #   ##   #
 X"1cce00", --     ###  ##  ###
 X"0edc00", --      ### ## ###
 X"03f000", --        ######
 X"00c000", --          ##
 X"03f000", --        ######
 X"0ffc00", --      ##########
 X"1cce00", --     ###  ##  ###
 X"08c400", --      #   ##   #
 X"00c000", --          ##
 X"00c000", --          ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 43 0x2B Plus sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"3fff80", --    ###############
 X"3fff80", --    ###############
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 44 0x2C Comma
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01c000", --         ###
 X"03e000", --        #####
 X"03e000", --        #####
 X"03e000", --        #####
 X"01e000", --         ####
 X"01e000", --         ####
 X"01c000", --         ###
 X"03c000", --        ####
 X"1f0000", --     #####
 X"1c0000", --     ###
 X"000000", -- 
-- char code 45 0x2D Hyphen-minus
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0ff800", --      #########
 X"0ff800", --      #########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 46 0x2E Full stop
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01c000", --         ###
 X"03e000", --        #####
 X"03e000", --        #####
 X"03e000", --        #####
 X"01c000", --         ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 47 0x2F Slash
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000600", --               ##
 X"000e00", --              ###
 X"000c00", --              ##
 X"001c00", --             ###
 X"001c00", --             ###
 X"001800", --             ##
 X"003800", --            ###
 X"003000", --            ##
 X"007000", --           ###
 X"006000", --           ##
 X"00e000", --          ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"018000", --         ##
 X"038000", --        ###
 X"030000", --        ##
 X"070000", --       ###
 X"060000", --       ##
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0c0000", --      ##
 X"1c0000", --     ###
 X"180000", --     ##
 X"380000", --    ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 48 0x30 Digit Zero
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03e000", --        #####
 X"0ff800", --      #########
 X"1e3c00", --     ####   ####
 X"3c1e00", --    ####     ####
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"700f00", --   ###        ####
 X"703f00", --   ###      ######
 X"707700", --   ###     ### ###
 X"70e700", --   ###    ###  ###
 X"738700", --   ###  ###    ###
 X"770700", --   ### ###     ###
 X"7e0700", --   ######      ###
 X"780700", --   ####        ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"3c1e00", --    ####     ####
 X"1e3c00", --     ####   ####
 X"0ff800", --      #########
 X"03e000", --        #####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 49 0x31 Digit One
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00e000", --          ###
 X"03e000", --        #####
 X"0ee000", --      ### ###
 X"1ce000", --     ###  ###
 X"38e000", --    ###   ###
 X"10e000", --     #    ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"1fff00", --     #############
 X"1fff00", --     #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 50 0x32 Digit Two
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"07e000", --       ######
 X"1ff000", --     #########
 X"387800", --    ###    ####
 X"103c00", --     #      ####
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"003c00", --            ####
 X"003800", --            ###
 X"007800", --           ####
 X"00f000", --          ####
 X"01e000", --         ####
 X"03c000", --        ####
 X"078000", --       ####
 X"0f0000", --      ####
 X"0e0000", --      ###
 X"1c0000", --     ###
 X"3ffe00", --    #############
 X"3ffe00", --    #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 51 0x33 Digit Three
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"07f000", --       #######
 X"0ffc00", --      ##########
 X"081c00", --      #      ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"001c00", --             ###
 X"003c00", --            ####
 X"03f000", --        ######
 X"03fc00", --        ########
 X"001e00", --             ####
 X"000f00", --              ####
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000e00", --              ###
 X"001e00", --             ####
 X"1ff800", --     ##########
 X"1fe000", --     ########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 52 0x34 Digit Four
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"003c00", --            ####
 X"007c00", --           #####
 X"00fc00", --          ######
 X"00dc00", --          ## ###
 X"01dc00", --         ### ###
 X"039c00", --        ###  ###
 X"039c00", --        ###  ###
 X"071c00", --       ###   ###
 X"0e1c00", --      ###    ###
 X"0e1c00", --      ###    ###
 X"1c1c00", --     ###     ###
 X"181c00", --     ##      ###
 X"381c00", --    ###      ###
 X"701c00", --   ###       ###
 X"7fff80", --   ################
 X"7fff80", --   ################
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 53 0x35 Digit Five
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1ff000", --     #########
 X"1ffc00", --     ###########
 X"001e00", --             ####
 X"000f00", --              ####
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000e00", --              ###
 X"003c00", --            ####
 X"1ff800", --     ##########
 X"1fe000", --     ########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 54 0x36 Digit Six
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00fc00", --          ######
 X"03fc00", --        ########
 X"078000", --       ####
 X"0e0000", --      ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"180000", --     ##
 X"380000", --    ###
 X"3bf800", --    ### #######
 X"3ffc00", --    ############
 X"3c1e00", --    ####     ####
 X"380f00", --    ###       ####
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"1c0700", --     ###       ###
 X"1c0e00", --     ###      ###
 X"0e1e00", --      ###    ####
 X"0ffc00", --      ##########
 X"03f000", --        ######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 55 0x37 Digit Seven
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3fff00", --    ##############
 X"3fff00", --    ##############
 X"000700", --               ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"003800", --            ###
 X"003800", --            ###
 X"007000", --           ###
 X"007000", --           ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"038000", --        ###
 X"038000", --        ###
 X"078000", --       ####
 X"070000", --       ###
 X"0f0000", --      ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 56 0x38 Digit Eight
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f800", --        #######
 X"0ffe00", --      ###########
 X"1c0e00", --     ###      ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3c0f00", --    ####      ####
 X"1e0e00", --     ####     ###
 X"0f3c00", --      ####  ####
 X"07f800", --       ########
 X"07f800", --       ########
 X"0f3c00", --      ####  ####
 X"1c0e00", --     ###      ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"1e1e00", --     ####    ####
 X"0ffc00", --      ##########
 X"07f000", --       #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 57 0x39 Digit Nine
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f000", --        ######
 X"0ff800", --      #########
 X"1e1c00", --     ####    ###
 X"1c0e00", --     ###      ###
 X"380e00", --    ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3c0700", --    ####       ###
 X"1e0f00", --     ####     ####
 X"0fff00", --      ############
 X"07f700", --       ####### ###
 X"000700", --               ###
 X"000600", --               ##
 X"000e00", --              ###
 X"001e00", --             ####
 X"003c00", --            ####
 X"007800", --           ####
 X"1ff000", --     #########
 X"1f8000", --     ######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 58 0x3A Colon
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"018000", --         ##
 X"03c000", --        ####
 X"03c000", --        ####
 X"03c000", --        ####
 X"018000", --         ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"018000", --         ##
 X"03c000", --        ####
 X"03c000", --        ####
 X"03c000", --        ####
 X"018000", --         ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 59 0x3B Semicolon
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00c000", --          ##
 X"01e000", --         ####
 X"01e000", --         ####
 X"01e000", --         ####
 X"00c000", --          ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00e000", --          ###
 X"01f000", --         #####
 X"01f000", --         #####
 X"01f000", --         #####
 X"00f000", --          ####
 X"00f000", --          ####
 X"00e000", --          ###
 X"01e000", --         ####
 X"0f8000", --      #####
 X"0e0000", --      ###
 X"000000", -- 
-- char code 60 0x3C Less-than sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000800", --              #
 X"001c00", --             ###
 X"007800", --           ####
 X"00f000", --          ####
 X"01e000", --         ####
 X"03c000", --        ####
 X"078000", --       ####
 X"0f0000", --      ####
 X"1e0000", --     ####
 X"1e0000", --     ####
 X"0f0000", --      ####
 X"078000", --       ####
 X"03c000", --        ####
 X"01e000", --         ####
 X"00f000", --          ####
 X"007800", --           ####
 X"001c00", --             ###
 X"000800", --              #
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 61 0x3D Equal sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3ffe00", --    #############
 X"3ffe00", --    #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3ffe00", --    #############
 X"3ffe00", --    #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 62 0x3E Greater-than sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"080000", --      #
 X"1c0000", --     ###
 X"0f0000", --      ####
 X"078000", --       ####
 X"03c000", --        ####
 X"01e000", --         ####
 X"00f000", --          ####
 X"007800", --           ####
 X"003c00", --            ####
 X"003c00", --            ####
 X"007800", --           ####
 X"00f000", --          ####
 X"01e000", --         ####
 X"03c000", --        ####
 X"078000", --       ####
 X"0f0000", --      ####
 X"1c0000", --     ###
 X"080000", --      #
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 63 0x3F Question mark
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"078000", --       ####
 X"07f000", --       #######
 X"007800", --           ####
 X"003c00", --            ####
 X"001c00", --             ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"001c00", --             ###
 X"01fc00", --         #######
 X"01f000", --         #####
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"000000", -- 
 X"000000", -- 
 X"018000", --         ##
 X"03c000", --        ####
 X"03c000", --        ####
 X"018000", --         ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 64 0x40 At sign
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01f800", --         ######
 X"03fc00", --        ########
 X"0f0e00", --      ####    ###
 X"0c0700", --      ##       ###
 X"180300", --     ##         ##
 X"380300", --    ###         ##
 X"300180", --    ##           ##
 X"700180", --   ###           ##
 X"61f980", --   ##    ######  ##
 X"63f980", --   ##   #######  ##
 X"673980", --   ##  ###  ###  ##
 X"c73980", --  ##   ###  ###  ##
 X"c63180", --  ##   ##   ##   ##
 X"ce3180", --  ##  ###   ##   ##
 X"ce3180", --  ##  ###   ##   ##
 X"ce3180", --  ##  ###   ##   ##
 X"ce3100", --  ##  ###   ##   #
 X"ce7300", --  ##  ###  ###  ##
 X"ce7300", --  ##  ###  ###  ##
 X"c7fe00", --  ##   ##########
 X"c79c00", --  ##   ####  ###
 X"e00000", --  ###
 X"600000", --   ##
 X"600000", --   ##
 X"300000", --    ##
 X"3c1800", --    ####     ##
 X"1ff800", --     ##########
 X"07e000", --       ######
-- char code 65 0x41 Latin Capital letter A
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01e000", --         ####
 X"03e000", --        #####
 X"036000", --        ## ##
 X"077000", --       ### ###
 X"077000", --       ### ###
 X"063000", --       ##   ##
 X"0e3800", --      ###   ###
 X"0e3800", --      ###   ###
 X"0c1800", --      ##     ##
 X"1c1c00", --     ###     ###
 X"1c1c00", --     ###     ###
 X"180e00", --     ##       ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"7fff00", --   ###############
 X"7fff00", --   ###############
 X"700700", --   ###         ###
 X"e00380", --  ###           ###
 X"e00380", --  ###           ###
 X"e00380", --  ###           ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 66 0x42 Latin Capital letter B
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3fe000", --    #########
 X"3ff800", --    ###########
 X"383800", --    ###     ###
 X"381c00", --    ###      ###
 X"381c00", --    ###      ###
 X"381c00", --    ###      ###
 X"381c00", --    ###      ###
 X"383800", --    ###     ###
 X"387800", --    ###    ####
 X"3fe000", --    #########
 X"3ff800", --    ###########
 X"383c00", --    ###     ####
 X"381e00", --    ###      ####
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"381e00", --    ###      ####
 X"383c00", --    ###     ####
 X"3ff800", --    ###########
 X"3fe000", --    #########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 67 0x43 Latin Capital letter C
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01fe00", --         ########
 X"07ff00", --       ###########
 X"0f0100", --      ####       #
 X"1c0000", --     ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"700000", --   ###
 X"700000", --   ###
 X"700000", --   ###
 X"700000", --   ###
 X"700000", --   ###
 X"700000", --   ###
 X"700000", --   ###
 X"380000", --    ###
 X"380000", --    ###
 X"1c0000", --     ###
 X"1f0300", --     #####      ##
 X"07ff00", --       ###########
 X"01fc00", --         #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 68 0x44 Latin Capital letter D
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3fe000", --    #########
 X"3ff800", --    ###########
 X"381e00", --    ###      ####
 X"380e00", --    ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380e00", --    ###       ###
 X"383c00", --    ###     ####
 X"3ff800", --    ###########
 X"3fe000", --    #########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 69 0x45 Latin Capital letter E
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 70 0x46 Latin Capital letter F
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 71 0x47 Latin Capital letter G
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01fe00", --         ########
 X"07ff00", --       ###########
 X"0f0100", --      ####       #
 X"1e0000", --     ####
 X"3c0000", --    ####
 X"380000", --    ###
 X"380000", --    ###
 X"700000", --   ###
 X"700000", --   ###
 X"707f00", --   ###     #######
 X"707f00", --   ###     #######
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"1c0700", --     ###       ###
 X"1f0700", --     #####     ###
 X"07ff00", --       ###########
 X"01fc00", --         #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 72 0x48 Latin Capital letter H
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3fff00", --    ##############
 X"3fff00", --    ##############
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 73 0x49 Latin Capital letter I
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3ffe00", --    #############
 X"3ffe00", --    #############
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"3ffe00", --    #############
 X"3ffe00", --    #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 74 0x4A Latin Capital letter J
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ffc00", --     ###########
 X"1ffc00", --     ###########
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"001c00", --             ###
 X"103800", --     #      ###
 X"187800", --     ##    ####
 X"0ff000", --      ########
 X"07c000", --       #####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 75 0x4B Latin Capital letter K
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"380700", --    ###        ###
 X"380e00", --    ###       ###
 X"381c00", --    ###      ###
 X"383800", --    ###     ###
 X"387000", --    ###    ###
 X"386000", --    ###    ##
 X"38e000", --    ###   ###
 X"39c000", --    ###  ###
 X"3b8000", --    ### ###
 X"3f0000", --    ######
 X"3f0000", --    ######
 X"3b8000", --    ### ###
 X"39c000", --    ###  ###
 X"38e000", --    ###   ###
 X"387000", --    ###    ###
 X"387800", --    ###    ####
 X"383c00", --    ###     ####
 X"381c00", --    ###      ###
 X"380e00", --    ###       ###
 X"380700", --    ###        ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 76 0x4C Latin Capital letter L
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0e0000", --      ###
 X"0fff00", --      ############
 X"0fff00", --      ############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 77 0x4D Latin Capital letter M
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3c0f00", --    ####      ####
 X"3c0f00", --    ####      ####
 X"3e0f00", --    #####     ####
 X"361b00", --    ## ##    ## ##
 X"361b00", --    ## ##    ## ##
 X"361300", --    ## ##    #  ##
 X"333300", --    ##  ##  ##  ##
 X"333300", --    ##  ##  ##  ##
 X"332300", --    ##  ##  #   ##
 X"31e300", --    ##   ####   ##
 X"31e300", --    ##   ####   ##
 X"31c300", --    ##   ###    ##
 X"30c300", --    ##    ##    ##
 X"300300", --    ##          ##
 X"300300", --    ##          ##
 X"300380", --    ##          ###
 X"300380", --    ##          ###
 X"300380", --    ##          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 78 0x4E Latin Capital letter N
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3c0700", --    ####       ###
 X"3e0700", --    #####      ###
 X"3e0700", --    #####      ###
 X"3e0700", --    #####      ###
 X"3b0700", --    ### ##     ###
 X"3b0700", --    ### ##     ###
 X"3b8700", --    ### ###    ###
 X"398700", --    ###  ##    ###
 X"39c700", --    ###  ###   ###
 X"38c700", --    ###   ##   ###
 X"38c700", --    ###   ##   ###
 X"38e700", --    ###   ###  ###
 X"386700", --    ###    ##  ###
 X"387700", --    ###    ### ###
 X"383700", --    ###     ## ###
 X"383700", --    ###     ## ###
 X"381f00", --    ###      #####
 X"381f00", --    ###      #####
 X"381f00", --    ###      #####
 X"380f00", --    ###       ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 79 0x4F Latin Capital letter O
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f000", --        ######
 X"0ffc00", --      ##########
 X"1e1e00", --     ####    ####
 X"1c0f00", --     ###      ####
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3c0e00", --    ####      ###
 X"1e1e00", --     ####    ####
 X"0ffc00", --      ##########
 X"03f000", --        ######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 80 0x50 Latin Capital letter P
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3ff000", --    ##########
 X"3ffc00", --    ############
 X"381e00", --    ###      ####
 X"380e00", --    ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380e00", --    ###       ###
 X"381c00", --    ###      ###
 X"3ff800", --    ###########
 X"3fe000", --    #########
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 81 0x51 Latin Capital letter Q
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f000", --        ######
 X"0ffc00", --      ##########
 X"1e1e00", --     ####    ####
 X"1c0f00", --     ###      ####
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3c0e00", --    ####      ###
 X"1e1e00", --     ####    ####
 X"0ffc00", --      ##########
 X"03f000", --        ######
 X"00e000", --          ###
 X"00e000", --          ###
 X"007000", --           ###
 X"007880", --           ####   #
 X"003fc0", --            ########
 X"001f80", --             ######
-- char code 82 0x52 Latin Capital letter R
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ff000", --     #########
 X"1ffc00", --     ###########
 X"1c1c00", --     ###     ###
 X"1c0e00", --     ###      ###
 X"1c0e00", --     ###      ###
 X"1c0e00", --     ###      ###
 X"1c0e00", --     ###      ###
 X"1c1e00", --     ###     ####
 X"1c3c00", --     ###    ####
 X"1ff800", --     ##########
 X"1fe000", --     ########
 X"1c7000", --     ###   ###
 X"1c3800", --     ###    ###
 X"1c3c00", --     ###    ####
 X"1c1c00", --     ###     ###
 X"1c1e00", --     ###     ####
 X"1c0e00", --     ###      ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0380", --     ###        ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 83 0x53 Latin Capital letter S
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f800", --        #######
 X"0ffe00", --      ###########
 X"1e0600", --     ####      ##
 X"3c0000", --    ####
 X"380000", --    ###
 X"380000", --    ###
 X"3c0000", --    ####
 X"1e0000", --     ####
 X"1f8000", --     ######
 X"07f000", --       #######
 X"01fc00", --         #######
 X"003e00", --            #####
 X"000f00", --              ####
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000f00", --              ####
 X"301e00", --    ##       ####
 X"3ffc00", --    ############
 X"0ff000", --      ########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 84 0x54 Latin Capital letter T
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"7fff00", --   ###############
 X"7fff00", --   ###############
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 85 0x55 Latin Capital letter U
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"1c0e00", --     ###      ###
 X"1e1e00", --     ####    ####
 X"0ffc00", --      ##########
 X"03f000", --        ######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 86 0x56 Latin Capital letter V
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"7001c0", --   ###           ###
 X"7001c0", --   ###           ###
 X"7001c0", --   ###           ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"3c0380", --    ####        ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1e0600", --     ####      ##
 X"0e0e00", --      ###     ###
 X"0e0e00", --      ###     ###
 X"070c00", --       ###    ##
 X"071c00", --       ###   ###
 X"071c00", --       ###   ###
 X"039800", --        ###  ##
 X"03b800", --        ### ###
 X"03b800", --        ### ###
 X"01f000", --         #####
 X"01f000", --         #####
 X"01e000", --         ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 87 0x57 Latin Capital letter W
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"700380", --   ###          ###
 X"70c380", --   ###    ##    ###
 X"70e380", --   ###    ###   ###
 X"71e380", --   ###   ####   ###
 X"31e300", --    ##   ####   ##
 X"31f300", --    ##   #####  ##
 X"333300", --    ##  ##  ##  ##
 X"333300", --    ##  ##  ##  ##
 X"333b00", --    ##  ##  ### ##
 X"3e1b00", --    #####    ## ##
 X"3e1b00", --    #####    ## ##
 X"3e1f00", --    #####    #####
 X"3c0f00", --    ####      ####
 X"3c0f00", --    ####      ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 88 0x58 Latin Capital letter X
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"780780", --   ####        ####
 X"380700", --    ###        ###
 X"1c0e00", --     ###      ###
 X"1e1e00", --     ####    ####
 X"0f1c00", --      ####   ###
 X"073800", --       ###  ###
 X"07f800", --       ########
 X"03f000", --        ######
 X"01e000", --         ####
 X"01e000", --         ####
 X"01f000", --         #####
 X"03f000", --        ######
 X"07f800", --       ########
 X"0f3c00", --      ####  ####
 X"0e1c00", --      ###    ###
 X"1e1e00", --     ####    ####
 X"3c0f00", --    ####      ####
 X"380700", --    ###        ###
 X"700780", --   ###         ####
 X"f003c0", --  ####          ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 89 0x59 Latin Capital letter Y
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"7001c0", --   ###           ###
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"0e0e00", --      ###     ###
 X"0f0e00", --      ####    ###
 X"071c00", --       ###   ###
 X"039800", --        ###  ##
 X"03b800", --        ### ###
 X"01f000", --         #####
 X"01f000", --         #####
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 90 0x5A Latin Capital letter Z
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3fff00", --    ##############
 X"3fff00", --    ##############
 X"000e00", --              ###
 X"000e00", --              ###
 X"001c00", --             ###
 X"003800", --            ###
 X"003800", --            ###
 X"007000", --           ###
 X"006000", --           ##
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"038000", --        ###
 X"070000", --       ###
 X"070000", --       ###
 X"0e0000", --      ###
 X"0c0000", --      ##
 X"1c0000", --     ###
 X"3fff00", --    ##############
 X"3fff00", --    ##############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 91 0x5B Left Square Bracket
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"07f800", --       ########
 X"07f800", --       ########
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"07f800", --       ########
 X"07f800", --       ########
-- char code 92 0x5C Backslash
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c0000", --     ###
 X"0c0000", --      ##
 X"0e0000", --      ###
 X"060000", --       ##
 X"070000", --       ###
 X"070000", --       ###
 X"030000", --        ##
 X"038000", --        ###
 X"018000", --         ##
 X"01c000", --         ###
 X"00c000", --          ##
 X"00e000", --          ###
 X"00e000", --          ###
 X"007000", --           ###
 X"007000", --           ###
 X"003000", --            ##
 X"003800", --            ###
 X"001800", --             ##
 X"001c00", --             ###
 X"000c00", --              ##
 X"000e00", --              ###
 X"000e00", --              ###
 X"000600", --               ##
 X"000700", --               ###
 X"000300", --                ##
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 93 0x5D Right Square Bracket
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"07f800", --       ########
 X"07f800", --       ########
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"07f800", --       ########
 X"07f800", --       ########
-- char code 94 0x5E Circumflex accent
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01c000", --         ###
 X"01e000", --         ####
 X"036000", --        ## ##
 X"077000", --       ### ###
 X"063000", --       ##   ##
 X"0e3800", --      ###   ###
 X"0c1800", --      ##     ##
 X"1c1c00", --     ###     ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 95 0x5F Low line
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"ffffc0", --  ##################
 X"ffffc0", --  ##################
-- char code 96 0x60 Grave accent
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0f0000", --      ####
 X"078000", --       ####
 X"03c000", --        ####
 X"01e000", --         ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 97 0x61 Latin Small Letter A
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"07f000", --       #######
 X"1ffc00", --     ###########
 X"181c00", --     ##      ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"000e00", --              ###
 X"07fe00", --       ##########
 X"1ffe00", --     ############
 X"1c0e00", --     ###      ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"381e00", --    ###      ####
 X"3c7e00", --    ####   ######
 X"1ffe00", --     ############
 X"0fce00", --      ######  ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 98 0x62 Latin Small Letter B
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c7c00", --     ###   #####
 X"1dfe00", --     ### ########
 X"1f8f00", --     ######   ####
 X"1f0700", --     #####     ###
 X"1e0380", --     ####       ###
 X"1c0380", --     ###        ###
 X"1c0380", --     ###        ###
 X"1c0380", --     ###        ###
 X"1c0380", --     ###        ###
 X"1c0380", --     ###        ###
 X"1c0380", --     ###        ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1e1e00", --     ####    ####
 X"1ffc00", --     ###########
 X"07f000", --       #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 99 0x63 Latin Small Letter C
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01f800", --         ######
 X"07fc00", --       #########
 X"0f0400", --      ####     #
 X"1e0000", --     ####
 X"1c0000", --     ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"3c0000", --    ####
 X"1c0000", --     ###
 X"0f0400", --      ####     #
 X"07fc00", --       #########
 X"03f800", --        #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 100 0x64 Latin Small Letter D
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"01ff00", --         #########
 X"07ff00", --       ###########
 X"0f0700", --      ####     ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380f00", --    ###       ####
 X"1c1f00", --     ###     #####
 X"1e3f00", --     ####   ######
 X"0ff700", --      ######## ###
 X"07c700", --       #####   ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 101 0x65 Latin Small Letter E
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f000", --        ######
 X"07fc00", --       #########
 X"0e1e00", --      ###    ####
 X"1c0e00", --     ###      ###
 X"1c0700", --     ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"3fff00", --    ##############
 X"3fff00", --    ##############
 X"380000", --    ###
 X"380000", --    ###
 X"380000", --    ###
 X"1c0000", --     ###
 X"1e0200", --     ####       #
 X"0ffe00", --      ###########
 X"03f800", --        #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 102 0x66 Latin Small Letter F
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"003f80", --            #######
 X"00ff80", --          #########
 X"01e000", --         ####
 X"03c000", --        ####
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"7fff00", --   ###############
 X"7fff00", --   ###############
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"038000", --        ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 103 0x67 Latin Small Letter G
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03ff80", --        ###########
 X"0fff80", --      #############
 X"1e3c00", --     ####   ####
 X"3c1e00", --    ####     ####
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"3c1e00", --    ####     ####
 X"1e3c00", --     ####   ####
 X"1ff800", --     ##########
 X"3be000", --    ### #####
 X"380000", --    ###
 X"380000", --    ###
 X"3c0000", --    ####
 X"1ffc00", --     ###########
 X"1ffe00", --     ############
 X"380f00", --    ###       ####
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"780e00", --   ####       ###
 X"3ffc00", --    ############
 X"0ff000", --      ########
-- char code 104 0x68 Latin Small Letter H
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c7800", --     ###   ####
 X"1dfe00", --     ### ########
 X"1f8e00", --     ######   ###
 X"1f0700", --     #####     ###
 X"1e0700", --     ####      ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 105 0x69 Latin Small Letter I
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"00c000", --          ##
 X"01e000", --         ####
 X"01e000", --         ####
 X"00c000", --          ##
 X"000000", -- 
 X"000000", -- 
 X"0fe000", --      #######
 X"0fe000", --      #######
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"1fff00", --     #############
 X"1fff00", --     #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 106 0x6A Latin Small Letter J
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"001800", --             ##
 X"003c00", --            ####
 X"003c00", --            ####
 X"001800", --             ##
 X"000000", -- 
 X"000000", -- 
 X"1ff800", --     ##########
 X"1ff800", --     ##########
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"003800", --            ###
 X"007000", --           ###
 X"20f000", --    #     ####
 X"3fe000", --    #########
 X"1f8000", --     ######
-- char code 107 0x6B Latin Small Letter K
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0700", --     ###       ###
 X"1c0e00", --     ###      ###
 X"1c1c00", --     ###     ###
 X"1c3800", --     ###    ###
 X"1c7000", --     ###   ###
 X"1ce000", --     ###  ###
 X"1dc000", --     ### ###
 X"1f8000", --     ######
 X"1dc000", --     ### ###
 X"1ce000", --     ###  ###
 X"1cf000", --     ###  ####
 X"1c7800", --     ###   ####
 X"1c3c00", --     ###    ####
 X"1c1e00", --     ###     ####
 X"1c0f00", --     ###      ####
 X"1c0780", --     ###       ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 108 0x6C Latin Small Letter L
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0fe000", --      #######
 X"0fe000", --      #######
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"1fff00", --     #############
 X"1fff00", --     #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 109 0x6D Latin Small Letter M
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"3bcf00", --    ### ####  ####
 X"3fdf00", --    ######## #####
 X"3cf380", --    ####  ####  ###
 X"3cf380", --    ####  ####  ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"38e380", --    ###   ###   ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 110 0x6E Latin Small Letter N
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c7c00", --     ###   #####
 X"1dfe00", --     ### ########
 X"1f8e00", --     ######   ###
 X"1f0700", --     #####     ###
 X"1e0700", --     ####      ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 111 0x6F Latin Small Letter O
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f000", --        ######
 X"0ff800", --      #########
 X"1c1c00", --     ###     ###
 X"380e00", --    ###       ###
 X"380f00", --    ###       ####
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"700700", --   ###         ###
 X"380e00", --    ###       ###
 X"380e00", --    ###       ###
 X"1c1c00", --     ###     ###
 X"0ff800", --      #########
 X"07e000", --       ######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 112 0x70 Latin Small Letter P
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1cf800", --     ###  #####
 X"1dfc00", --     ### #######
 X"1f8e00", --     ######   ###
 X"1e0e00", --     ####     ###
 X"1e0700", --     ####      ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0e00", --     ###      ###
 X"1c0e00", --     ###      ###
 X"1c1c00", --     ###     ###
 X"1ff800", --     ##########
 X"1ff000", --     #########
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
-- char code 113 0x71 Latin Small Letter Q
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"01ff00", --         #########
 X"07ff00", --       ###########
 X"0f0700", --      ####     ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380700", --    ###        ###
 X"380f00", --    ###       ####
 X"1c1f00", --     ###     #####
 X"1e3f00", --     ####   ######
 X"0ff700", --      ######## ###
 X"07c700", --       #####   ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
 X"000700", --               ###
-- char code 114 0x72 Latin Small Letter R
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c7c00", --     ###   #####
 X"1dfe00", --     ### ########
 X"1f8e00", --     ######   ###
 X"1f0700", --     #####     ###
 X"1e0700", --     ####      ###
 X"1c0700", --     ###       ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 115 0x73 Latin Small Letter S
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"03f800", --        #######
 X"0ffc00", --      ##########
 X"0e0400", --      ###      #
 X"1c0000", --     ###
 X"1c0000", --     ###
 X"1e0000", --     ####
 X"0f8000", --      #####
 X"07f000", --       #######
 X"03fc00", --        ########
 X"003e00", --            #####
 X"001e00", --             ####
 X"000e00", --              ###
 X"000e00", --              ###
 X"181c00", --     ##      ###
 X"1ffc00", --     ###########
 X"0ff000", --      ########
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 116 0x74 Latin Small Letter T
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"030000", --        ##
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"7ffe00", --   ##############
 X"7ffe00", --   ##############
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"070000", --       ###
 X"038000", --        ###
 X"03c000", --        ####
 X"01fe00", --         ########
 X"00fe00", --          #######
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 117 0x75 Latin Small Letter U
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"1c0f00", --     ###      ####
 X"1c1f00", --     ###     #####
 X"0e3f00", --      ###   ######
 X"0ff700", --      ######## ###
 X"07c700", --       #####   ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 118 0x76 Latin Small Letter V
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"380300", --    ###         ##
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"0e0e00", --      ###     ###
 X"0e0e00", --      ###     ###
 X"0e0c00", --      ###     ##
 X"071c00", --       ###   ###
 X"071c00", --       ###   ###
 X"031800", --        ##   ##
 X"03b800", --        ### ###
 X"03b000", --        ### ##
 X"01b000", --         ## ##
 X"01f000", --         #####
 X"00e000", --          ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 119 0x77 Latin Small Letter W
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"600300", --   ##           ##
 X"600300", --   ##           ##
 X"600300", --   ##           ##
 X"600700", --   ##          ###
 X"71c700", --   ###   ###   ###
 X"71c700", --   ###   ###   ###
 X"71c700", --   ###   ###   ###
 X"736600", --   ###  ## ##  ##
 X"336600", --    ##  ## ##  ##
 X"336600", --    ##  ## ##  ##
 X"326600", --    ##  #  ##  ##
 X"363600", --    ## ##   ## ##
 X"363600", --    ## ##   ## ##
 X"3e3e00", --    #####   #####
 X"3c1e00", --    ####     ####
 X"3c1c00", --    ####     ###
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 120 0x78 Latin Small Letter X
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"780f00", --   ####       ####
 X"3c0e00", --    ####      ###
 X"1c1c00", --     ###     ###
 X"0e3800", --      ###   ###
 X"0f3800", --      ####  ###
 X"077000", --       ### ###
 X"03e000", --        #####
 X"01e000", --         ####
 X"03e000", --        #####
 X"03f000", --        ######
 X"077800", --       ### ####
 X"0e3800", --      ###   ###
 X"0e1c00", --      ###    ###
 X"1c0e00", --     ###      ###
 X"3c0f00", --    ####      ####
 X"780780", --   ####        ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 121 0x79 Latin Small Letter Y
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"380380", --    ###         ###
 X"380380", --    ###         ###
 X"1c0300", --     ###        ##
 X"1c0700", --     ###       ###
 X"1c0700", --     ###       ###
 X"0e0e00", --      ###     ###
 X"0e0e00", --      ###     ###
 X"060c00", --       ##     ##
 X"071c00", --       ###   ###
 X"071800", --       ###   ##
 X"031800", --        ##   ##
 X"03b000", --        ### ##
 X"01b000", --         ## ##
 X"01f000", --         #####
 X"01e000", --         ####
 X"00e000", --          ###
 X"00c000", --          ##
 X"01c000", --         ###
 X"038000", --        ###
 X"070000", --       ###
 X"7f0000", --   #######
 X"7c0000", --   #####
-- char code 122 0x7A Latin Small Letter Z
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1ffe00", --     ############
 X"1ffe00", --     ############
 X"001c00", --             ###
 X"001c00", --             ###
 X"003800", --            ###
 X"007000", --           ###
 X"007000", --           ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"018000", --         ##
 X"038000", --        ###
 X"070000", --       ###
 X"060000", --       ##
 X"0e0000", --      ###
 X"1fff00", --     #############
 X"1fff00", --     #############
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 123 0x7B Left Curly Bracket
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"003c00", --            ####
 X"00fc00", --          ######
 X"00e000", --          ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"038000", --        ###
 X"1f0000", --     #####
 X"1f0000", --     #####
 X"038000", --        ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"01c000", --         ###
 X"00e000", --          ###
 X"00fc00", --          ######
 X"003c00", --            ####
-- char code 124 0x7C Vertical bar
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
-- char code 125 0x7D Right Curly Bracket
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"0f0000", --      ####
 X"0fc000", --      ######
 X"01c000", --         ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"007000", --           ###
 X"003e00", --            #####
 X"003e00", --            #####
 X"007000", --           ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"00e000", --          ###
 X"01c000", --         ###
 X"0fc000", --      ######
 X"0f0000", --      ####
-- char code 126 0x7E Tilde
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"1e0000", --     ####
 X"3f8380", --    #######     ###
 X"79c380", --   ####  ###    ###
 X"70e780", --   ###    ###  ####
 X"707f00", --   ###     #######
 X"001e00", --             ####
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
 X"000000", -- 
-- char code 127 0x7F Delete
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 
 X"000000",  -- 

 X"000000",  -- 
 X"000000",  -- 
 X"000000",  --  
 X"000000"   --  
 );
begin
-- Do not change the process!!! It has the structure that converts to M9k memory blocks
pixelOn: process (clk)
    variable ix:integer range 0 to ROM'LENGTH-1;
	begin
		ix:=to_integer(unsigned(addr));
		if rising_edge(clk) then
			-- Read from Rom
			fontRow <= ROM(ix);
		end if;
	end process;
	
end Behavioral;