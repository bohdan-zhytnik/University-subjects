library verilog;
use verilog.vl_types.all;
entity MorseBDF_prototype_vlg_vec_tst is
end MorseBDF_prototype_vlg_vec_tst;
