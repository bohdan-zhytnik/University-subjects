library verilog;
use verilog.vl_types.all;
entity majorita3_vlg_vec_tst is
end majorita3_vlg_vec_tst;
