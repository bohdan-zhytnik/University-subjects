library verilog;
use verilog.vl_types.all;
entity MorseBDF_vlg_vec_tst is
end MorseBDF_vlg_vec_tst;
