library verilog;
use verilog.vl_types.all;
entity majorita3n_vlg_vec_tst is
end majorita3n_vlg_vec_tst;
